module SHA3(
    in, more, input_valid, out, next, ready
);
input [1087:0] in;
input more, input_valid,;
output [255:0] out;
output next, ready;

Ffunction keccak_f(

);

//comb
always @() begin
    
end

//seq
always @(posedge clk) begin
    
end

endmodule